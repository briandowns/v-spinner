module spinner

import os
import sync
import term
import time

// spinner maintains the state for the spinner.
@[noinit]
struct Spinner {
mut:
	mu                sync.Mutex
	char_set          []string
	delay             time.Duration
	prefix            string
	suffix            string
	final_message     string
	last_output_plain string
	stop_chan         chan bool
	active            bool
	hide_cursor       bool
}

// Spinner.new creates a new value with the given
// character set.
pub fn Spinner.new(char_set int) Spinner {
	mut mu := sync.new_mutex()
	mu.init()

	return Spinner{
		mu: mu
		char_set: character_sets[char_set].clone()
		delay: 100 * time.millisecond
		hide_cursor: false
		active: false
	}
}

// set_hide_cursor sets the given value to hide or
// not hide the cursor.
pub fn (mut s Spinner) set_hide_cursor(hide bool) {
	s.mu.@lock()
	s.hide_cursor = hide
	s.mu.unlock()
}

// set_delay sets the delay to the given value.
pub fn (mut s Spinner) set_delay(delay time.Duration) {
	s.mu.@lock()
	s.delay = delay
	s.mu.unlock()
}

// set_prefix sets the prefix field with
// the given value.
pub fn (mut s Spinner) set_prefix(prefix string) {
	s.mu.@lock()
	s.prefix = prefix
	s.mu.unlock()
}

// set_suffix sets the suffix field with
// the given value.
pub fn (mut s Spinner) set_suffix(suffix string) {
	s.mu.@lock()
	s.suffix = suffix
	s.mu.unlock()
}

// set_final_message sets the final message field with
// the given value.
pub fn (mut s Spinner) set_final_message(fm string) {
	s.mu.@lock()
	s.final_message = fm
	s.mu.unlock()
}

// set_char_set sets the character set field with
// the given value.
pub fn (mut s Spinner) set_char_set(cs int) {
	s.mu.@lock()
	s.char_set = character_sets[cs].close()
	s.mu.unlock()
}

// start starts the spinner.
pub fn (mut s Spinner) start() {
	s.mu.@lock()

	if s.active || os.is_atty(os.stdout().fd) != 1 {
		s.mu.unlock()
		return
	}

	if s.hide_cursor {
		term.hide_cursor()
	}

	s.active = true
	s.mu.unlock()

	spawn fn (s Spinner) {
		for {
			for c in s.char_set {
				select {
					_ := <-s.stop_chan {
						return
					}
					10 * time.millisecond {
						print('\r${s.prefix}${c}${s.suffix}')
						os.flush()
						time.sleep(s.delay)
					}
				}
			}
		}

		print('\n')
	}(s)
}

// stop stops the spinner.
pub fn (mut s Spinner) stop() {
	s.mu.@lock()
	defer {
		s.mu.unlock()
	}

	if s.active {
		s.active = false
		// stop the spinner

		if s.hide_cursor {
			term.show_cursor()
		}

		s.erase()

		if s.final_message != '' {
			print('\r' + s.final_message)
		}
	}
}

// restart
pub fn (mut s Spinner) restart() {
	s.stop()
	s.start()
}

pub fn (mut s Spinner) reverse() {
	s.mu.@lock()
	s.char_set.reverse_in_place()
	s.mu.unlock()
}

// erase
fn (mut s Spinner) erase() {
	print('\r')
}

// fn main() {
// 	mut s := Spinner.new(35)
// 	s.set_hide_cursor(true)
// 	s.start()
// 	time.sleep(10 * time.second) // fake some work
// 	s.stop()

// 	println('we stopped the spinner!')
// }

const character_sets = {
	0:  ['←', '↖', '↑', '↗', '→', '↘', '↓', '↙']
	1:  ['▁', '▃', '▄', '▅', '▆', '▇', '█', '▇', '▆', '▅', '▄', '▃', '▁']
	2:  ['▖', '▘', '▝', '▗']
	3:  ['┤', '┘', '┴', '└', '├', '┌', '┬', '┐']
	4:  ['◢', '◣', '◤', '◥']
	5:  ['◰', '◳', '◲', '◱']
	6:  ['◴', '◷', '◶', '◵']
	7:  ['◐', '◓', '◑', '◒']
	8:  ['.', 'o', 'O', '@', '*']
	9:  ['|', '/', '-', '\\']
	10: ['◡◡', '⊙⊙', '◠◠']
	11: ['⣾', '⣽', '⣻', '⢿', '⡿', '⣟', '⣯', '⣷']
	12: [">))'>", " >))'>", "  >))'>", "   >))'>", "    >))'>", "   <'((<", "  <'((<", " <'((<"]
	13: ['⠁', '⠂', '⠄', '⡀', '⢀', '⠠', '⠐', '⠈']
	14: ['⠋', '⠙', '⠹', '⠸', '⠼', '⠴', '⠦', '⠧', '⠇', '⠏']
	15: ['a', 'b', 'c', 'd', 'e', 'f', 'g', 'h', 'i', 'j', 'k', 'l', 'm', 'n', 'o', 'p', 'q', 'r',
		's', 't', 'u', 'v', 'w', 'x', 'y', 'z']
	16: ['▉', '▊', '▋', '▌', '▍', '▎', '▏', '▎', '▍', '▌', '▋', '▊', '▉']
	17: ['■', '□', '▪', '▫']
	18: ['←', '↑', '→', '↓']
	19: ['╫', '╪']
	20: ['⇐', '⇖', '⇑', '⇗', '⇒', '⇘', '⇓', '⇙']
	21: ['⠁', '⠁', '⠉', '⠙', '⠚', '⠒', '⠂', '⠂', '⠒', '⠲', '⠴', '⠤', '⠄',
		'⠄', '⠤', '⠠', '⠠', '⠤', '⠦', '⠖', '⠒', '⠐', '⠐', '⠒', '⠓', '⠋',
		'⠉', '⠈', '⠈']
	22: ['⠈', '⠉', '⠋', '⠓', '⠒', '⠐', '⠐', '⠒', '⠖', '⠦', '⠤', '⠠', '⠠',
		'⠤', '⠦', '⠖', '⠒', '⠐', '⠐', '⠒', '⠓', '⠋', '⠉', '⠈']
	23: ['⠁', '⠉', '⠙', '⠚', '⠒', '⠂', '⠂', '⠒', '⠲', '⠴', '⠤', '⠄', '⠄',
		'⠤', '⠴', '⠲', '⠒', '⠂', '⠂', '⠒', '⠚', '⠙', '⠉', '⠁']
	24: ['⠋', '⠙', '⠚', '⠒', '⠂', '⠂', '⠒', '⠲', '⠴', '⠦', '⠖', '⠒', '⠐',
		'⠐', '⠒', '⠓', '⠋']
	25: ['ｦ', 'ｧ', 'ｨ', 'ｩ', 'ｪ', 'ｫ', 'ｬ', 'ｭ', 'ｮ', 'ｯ', 'ｱ', 'ｲ', 'ｳ',
		'ｴ', 'ｵ', 'ｶ', 'ｷ', 'ｸ', 'ｹ', 'ｺ', 'ｻ', 'ｼ', 'ｽ', 'ｾ', 'ｿ', 'ﾀ',
		'ﾁ', 'ﾂ', 'ﾃ', 'ﾄ', 'ﾅ', 'ﾆ', 'ﾇ', 'ﾈ', 'ﾉ', 'ﾊ', 'ﾋ', 'ﾌ', 'ﾍ',
		'ﾎ', 'ﾏ', 'ﾐ', 'ﾑ', 'ﾒ', 'ﾓ', 'ﾔ', 'ﾕ', 'ﾖ', 'ﾗ', 'ﾘ', 'ﾙ', 'ﾚ',
		'ﾛ', 'ﾜ', 'ﾝ']
	26: ['.', '..', '...']
	27: ['▁', '▂', '▃', '▄', '▅', '▆', '▇', '█', '▉', '▊', '▋', '▌', '▍',
		'▎', '▏', '▏', '▎', '▍', '▌', '▋', '▊', '▉', '█', '▇', '▆', '▅',
		'▄', '▃', '▂', '▁']
	28: ['.', 'o', 'O', '°', 'O', 'o', '.']
	29: ['+', 'x']
	30: ['v', '<', '^', '>']
	31: ['>>--->', ' >>--->', '  >>--->', '   >>--->', '    >>--->', '    <---<<', '   <---<<',
		'  <---<<', ' <---<<', '<---<<']
	32: ['|', '||', '|||', '||||', '|||||', '|||||||', '||||||||', '|||||||', '||||||', '|||||',
		'||||', '|||', '||', '|']
	33: ['[          ]', '[=         ]', '[==        ]', '[===       ]', '[====      ]',
		'[=====     ]', '[======    ]', '[=======   ]', '[========  ]', '[========= ]',
		'[==========]']
	34: ['(*---------)', '(-*--------)', '(--*-------)', '(---*------)', '(----*-----)',
		'(-----*----)', '(------*---)', '(-------*--)', '(--------*-)', '(---------*)']
	35: ['█▒▒▒▒▒▒▒▒▒', '███▒▒▒▒▒▒▒',
		'█████▒▒▒▒▒', '███████▒▒▒',
		'██████████']
	36: ['[                    ]', '[=>                  ]', '[===>                ]',
		'[=====>              ]', '[======>             ]', '[========>           ]',
		'[==========>         ]', '[============>       ]', '[==============>     ]',
		'[================>   ]', '[==================> ]', '[===================>]']
	39: ['🌍', '🌎', '🌏']
	40: ['◜', '◝', '◞', '◟']
	41: ['⬒', '⬔', '⬓', '⬕']
	42: ['⬖', '⬘', '⬗', '⬙']
	43: ['[>>>          >]', '[]>>>>        []', '[]  >>>>      []', '[]    >>>>    []',
		'[]      >>>>  []', '[]        >>>>[]', '[>>          >>]']
	44: ['♠', '♣', '♥', '♦']
	45: ['➞', '➟', '➠', '➡', '➠', '➟']
	46: ['  |  ', ' \\   ', '_    ', ' \\   ', '  |  ', '   / ', '    _', '   / ']
	47: ['  . . . .', '.   . . .', '. .   . .', '. . .   .', '. . . .  ', '. . . . .']
	48: [' |     ', '  /    ', '   _   ', '    \\  ', '     | ', '    \\  ', '   _   ', '  /    ']
	49: ['⎺', '⎻', '⎼', '⎽', '⎼', '⎻']
	50: ['▹▹▹▹▹', '▸▹▹▹▹', '▹▸▹▹▹', '▹▹▸▹▹',
		'▹▹▹▸▹', '▹▹▹▹▸']
	51: ['[    ]', '[   =]', '[  ==]', '[ ===]', '[====]', '[=== ]', '[==  ]', '[=   ]']
	52: ['( ●    )', '(  ●   )', '(   ●  )', '(    ● )', '(     ●)', '(    ● )',
		'(   ●  )', '(  ●   )', '( ●    )']
	53: ['✶', '✸', '✹', '✺', '✹', '✷']
	54: ['▐|\\____________▌', '▐_|\\___________▌', '▐__|\\__________▌',
		'▐___|\\_________▌', '▐____|\\________▌', '▐_____|\\_______▌',
		'▐______|\\______▌', '▐_______|\\_____▌', '▐________|\\____▌',
		'▐_________|\\___▌', '▐__________|\\__▌', '▐___________|\\_▌',
		'▐____________|\\▌', '▐____________/|▌', '▐___________/|_▌',
		'▐__________/|__▌', '▐_________/|___▌', '▐________/|____▌',
		'▐_______/|_____▌', '▐______/|______▌', '▐_____/|_______▌',
		'▐____/|________▌', '▐___/|_________▌', '▐__/|__________▌',
		'▐_/|___________▌', '▐/|____________▌']
	55: ['▐⠂       ▌', '▐⠈       ▌', '▐ ⠂      ▌', '▐ ⠠      ▌',
		'▐  ⡀     ▌', '▐  ⠠     ▌', '▐   ⠂    ▌', '▐   ⠈    ▌',
		'▐    ⠂   ▌', '▐    ⠠   ▌', '▐     ⡀  ▌', '▐     ⠠  ▌',
		'▐      ⠂ ▌', '▐      ⠈ ▌', '▐       ⠂▌', '▐       ⠠▌',
		'▐       ⡀▌', '▐      ⠠ ▌', '▐      ⠂ ▌', '▐     ⠈  ▌',
		'▐     ⠂  ▌', '▐    ⠠   ▌', '▐    ⡀   ▌', '▐   ⠠    ▌',
		'▐   ⠂    ▌', '▐  ⠈     ▌', '▐  ⠂     ▌', '▐ ⠠      ▌',
		'▐ ⡀      ▌', '▐⠠       ▌']
	56: ['¿', '?']
	57: ['⢹', '⢺', '⢼', '⣸', '⣇', '⡧', '⡗', '⡏']
	58: ['⢄', '⢂', '⢁', '⡁', '⡈', '⡐', '⡠']
	59: ['.  ', '.. ', '...', ' ..', '  .', '   ']
	60: ['.', 'o', 'O', '°', 'O', 'o', '.']
	61: ['▓', '▒', '░']
	62: ['▌', '▀', '▐', '▄']
	63: ['⊶', '⊷']
	64: ['▪', '▫']
	65: ['□', '■']
	66: ['▮', '▯']
	67: ['-', '=', '≡']
	68: ['d', 'q', 'p', 'b']
	69: ['∙∙∙', '●∙∙', '∙●∙', '∙∙●', '∙∙∙']
	70: ['🌑 ', '🌒 ', '🌓 ', '🌔 ', '🌕 ', '🌖 ', '🌗 ', '🌘 ']
	71: ['☗', '☖']
	72: ['⧇', '⧆']
	73: ['◉', '◎']
	74: ['㊂', '㊀', '㊁']
	75: ['⦾', '⦿']
	76: ['ဝ', '၀']
	77: ['▌', '▀', '▐▄']
	78: ['⠈⠁', '⠈⠑', '⠈⠱', '⠈⡱', '⢀⡱', '⢄⡱', '⢄⡱', '⢆⡱', '⢎⡱',
		'⢎⡰', '⢎⡠', '⢎⡀', '⢎⠁', '⠎⠁', '⠊⠁']
	79: ['________', '-_______', '_-______', '__-_____', '___-____', '____-___', '_____-__',
		'______-_', '_______-', '________', '_______-', '______-_', '_____-__', '____-___',
		'___-____', '__-_____', '_-______', '-_______', '________']
	80: ['|_______', '_/______', '__-_____', '___\\____', '____|___', '_____/__', '______-_',
		'_______\\', '_______|', '______\\_', '_____-__', '____/___', '___|____', '__\\_____',
		'_-______']
	81: ['□', '◱', '◧', '▣', '■']
	82: ['□', '◱', '▨', '▩', '■']
	83: ['░', '▒', '▓', '█']
	84: ['░', '█']
	85: ['⚪', '⚫']
	86: ['◯', '⬤']
	87: ['▱', '▰']
	88: ['➊', '➋', '➌', '➍', '➎', '➏', '➐', '➑', '➒', '➓']
	89: ['½', '⅓', '⅔', '¼', '¾', '⅛', '⅜', '⅝', '⅞']
	90: ['↞', '↟', '↠', '↡']
}
